weaver@pslab01.slac.stanford.edu.80142:1513882908